`timescale 1ns / 1ps
///////////////////////////////////////////////////////////////////////////////
// Company:         HomeDL
// Engineer:        ko
//
// Create Date:     23:22:20 02/27/2026
// Design Name:     pong_p_chu
// Module Name:     e_4_7_7
// Project Name:    -
// Target Devices:  -
// Tool versions:   -
// Description:     Stack
//
// Dependencies:    -
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments: -
//
///////////////////////////////////////////////////////////////////////////////
module e_4_7_7 (data_out, data_in, clock, reset, push, pop);
output data_out;
input data_in, clock, reset, push, pop;

wire [7:0] data_out, data_in;
wire clock, reset, push, pop;

endmodule
