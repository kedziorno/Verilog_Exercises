`timescale 1ns / 1ps
///////////////////////////////////////////////////////////////////////////////
// Company:         HomeDL
// Engineer:        ko
//
// Create Date:     20:54:40 02/13/2026
// Design Name:     pong_p_chu
// Module Name:     e_4_7_4
// Project Name:    -
// Target Devices:  -
// Tool versions:   -
// Description:     Heartbeat circuit
//
// Dependencies:    -
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments: -
//
///////////////////////////////////////////////////////////////////////////////
module e_4_7_4 (anode, segment, clock, reset);
output anode, segment;
input clock, reset;

wire [3:0] anode;
wire [6:0] segment;
wire clock, reset;


endmodule
