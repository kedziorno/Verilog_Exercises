// Verilog test fixture created from schematic /home/user/_WORKSPACE_/kedziorno/pong_p_chu/sch_e_2_9_2_7.sch - Sat Jan 17 18:58:37 2026
// ko, HomeDL
// 4-to-16 decoder with enable

`timescale 1ns / 1ps

module tb_sch_e_2_9_2_7();

// Inputs
reg i0;
reg i1;
reg i3;
reg i2;
reg en;

// Output
wire o0;
wire o1;
wire o2;
wire o3;
wire o4;
wire o5;
wire o6;
wire o7;
wire o8;
wire o9;
wire o10;
wire o11;
wire o12;
wire o13;
wire o14;
wire o15;

// Bidirs

// Instantiate the UUT
sch_e_2_9_2_7 UUT (
.i0(i0), .i1(i1), .i3(i3), .i2(i2), 
.en(en), 
.o0(o0), .o1(o1), .o2(o2), .o3(o3), 
.o4(o4), .o5(o5), .o6(o6), .o7(o7), 
.o8(o8), .o9(o9), .o10(o10), .o11(o11), 
.o12(o12), .o13(o13), .o14(o14), .o15(o15));

// Initialize Inputs
initial begin
i0 = 0;
i1 = 0;
i3 = 0;
i2 = 0;
en = 0;
#100;

en = 1; i3 = 0; i2 = 0; i1 = 0; i0 = 0; #100;
en = 1; i3 = 0; i2 = 0; i1 = 0; i0 = 1; #100;
en = 1; i3 = 0; i2 = 0; i1 = 1; i0 = 0; #100;
en = 1; i3 = 0; i2 = 0; i1 = 1; i0 = 1; #100;
en = 1; i3 = 0; i2 = 1; i1 = 0; i0 = 0; #100;
en = 1; i3 = 0; i2 = 1; i1 = 0; i0 = 1; #100;
en = 1; i3 = 0; i2 = 1; i1 = 1; i0 = 0; #100;
en = 1; i3 = 0; i2 = 1; i1 = 1; i0 = 1; #100;
en = 1; i3 = 1; i2 = 0; i1 = 0; i0 = 0; #100;
en = 1; i3 = 1; i2 = 0; i1 = 0; i0 = 1; #100;
en = 1; i3 = 1; i2 = 0; i1 = 1; i0 = 0; #100;
en = 1; i3 = 1; i2 = 0; i1 = 1; i0 = 1; #100;
en = 1; i3 = 1; i2 = 1; i1 = 0; i0 = 0; #100;
en = 1; i3 = 1; i2 = 1; i1 = 0; i0 = 1; #100;
en = 1; i3 = 1; i2 = 1; i1 = 1; i0 = 0; #100;
en = 1; i3 = 1; i2 = 1; i1 = 1; i0 = 1; #100;

en = 0; i3 = 0; i2 = 0; i1 = 0; i0 = 0; #100;
en = 0; i3 = 0; i2 = 0; i1 = 0; i0 = 1; #100;
en = 0; i3 = 0; i2 = 0; i1 = 1; i0 = 0; #100;
en = 0; i3 = 0; i2 = 0; i1 = 1; i0 = 1; #100;
en = 0; i3 = 0; i2 = 1; i1 = 0; i0 = 0; #100;
en = 0; i3 = 0; i2 = 1; i1 = 0; i0 = 1; #100;
en = 0; i3 = 0; i2 = 1; i1 = 1; i0 = 0; #100;
en = 0; i3 = 0; i2 = 1; i1 = 1; i0 = 1; #100;
en = 0; i3 = 1; i2 = 0; i1 = 0; i0 = 0; #100;
en = 0; i3 = 1; i2 = 0; i1 = 0; i0 = 1; #100;
en = 0; i3 = 1; i2 = 0; i1 = 1; i0 = 0; #100;
en = 0; i3 = 1; i2 = 0; i1 = 1; i0 = 1; #100;
en = 0; i3 = 1; i2 = 1; i1 = 0; i0 = 0; #100;
en = 0; i3 = 1; i2 = 1; i1 = 0; i0 = 1; #100;
en = 0; i3 = 1; i2 = 1; i1 = 1; i0 = 0; #100;
en = 0; i3 = 1; i2 = 1; i1 = 1; i0 = 1; #100;

en = 1; i3 = 0; i2 = 0; i1 = 0; i0 = 0; #100;
en = 0; i3 = 0; i2 = 0; i1 = 0; i0 = 1; #100;
en = 1; i3 = 0; i2 = 0; i1 = 1; i0 = 0; #100;
en = 0; i3 = 0; i2 = 0; i1 = 1; i0 = 1; #100;
en = 1; i3 = 0; i2 = 1; i1 = 0; i0 = 0; #100;
en = 0; i3 = 0; i2 = 1; i1 = 0; i0 = 1; #100;
en = 1; i3 = 0; i2 = 1; i1 = 1; i0 = 0; #100;
en = 0; i3 = 0; i2 = 1; i1 = 1; i0 = 1; #100;
en = 1; i3 = 1; i2 = 0; i1 = 0; i0 = 0; #100;
en = 0; i3 = 1; i2 = 0; i1 = 0; i0 = 1; #100;
en = 1; i3 = 1; i2 = 0; i1 = 1; i0 = 0; #100;
en = 0; i3 = 1; i2 = 0; i1 = 1; i0 = 1; #100;
en = 1; i3 = 1; i2 = 1; i1 = 0; i0 = 0; #100;
en = 0; i3 = 1; i2 = 1; i1 = 0; i0 = 1; #100;
en = 1; i3 = 1; i2 = 1; i1 = 1; i0 = 0; #100;
en = 0; i3 = 1; i2 = 1; i1 = 1; i0 = 1; #100;

en = 0; i3 = 0; i2 = 0; i1 = 0; i0 = 0; #100;
en = 1; i3 = 0; i2 = 0; i1 = 0; i0 = 1; #100;
en = 0; i3 = 0; i2 = 0; i1 = 1; i0 = 0; #100;
en = 1; i3 = 0; i2 = 0; i1 = 1; i0 = 1; #100;
en = 0; i3 = 0; i2 = 1; i1 = 0; i0 = 0; #100;
en = 1; i3 = 0; i2 = 1; i1 = 0; i0 = 1; #100;
en = 0; i3 = 0; i2 = 1; i1 = 1; i0 = 0; #100;
en = 1; i3 = 0; i2 = 1; i1 = 1; i0 = 1; #100;
en = 0; i3 = 1; i2 = 0; i1 = 0; i0 = 0; #100;
en = 1; i3 = 1; i2 = 0; i1 = 0; i0 = 1; #100;
en = 0; i3 = 1; i2 = 0; i1 = 1; i0 = 0; #100;
en = 1; i3 = 1; i2 = 0; i1 = 1; i0 = 1; #100;
en = 0; i3 = 1; i2 = 1; i1 = 0; i0 = 0; #100;
en = 1; i3 = 1; i2 = 1; i1 = 0; i0 = 1; #100;
en = 0; i3 = 1; i2 = 1; i1 = 1; i0 = 0; #100;
en = 1; i3 = 1; i2 = 1; i1 = 1; i0 = 1; #100;

$finish;
end

endmodule
